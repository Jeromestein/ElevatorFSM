module LiftFSM (
    ports
);
    
    
endmodule